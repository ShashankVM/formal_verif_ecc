module error_inject #(DATA_WIDTH=39) (
 logic [DATA_WIDTH-1:0] din, logic error_pos1, output logic [DATA_WIDTH-1:0] dout
 );
